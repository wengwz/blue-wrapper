typedef 8 AXI4_LEN_WIDTH;
typedef 3 AXI4_SIZE_WIDTH;
typedef 2 AXI4_BURST_WIDTH;
typedef 1 AXI4_LOCK_WIDTH;
typedef 4 AXI4_CACHE_WIDTH;
typedef 3 AXI4_PROT_WIDTH;
typedef 4 AXI4_QOS_WIDTH;
typedef 2 AXI4_RESP_WIDTH;

typedef 8 BYTE_WIDTH;